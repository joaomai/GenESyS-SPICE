.model diode D (Is=1E-16 vj=0.7)
