GenESyS generated circuit

.include ./diode.cir

Vs1 net_1 gnd sin(0 12.000000 60.000000 ) 
D1 net_2 net_1 diode 
D2 net_2 gnd diode 
D3 net_1 net_3 diode 
D4 gnd net_2 diode 
C1 net_3 net_2 9.999999m  
R1 net_3 net_2 1.000000K  

.control
tran 1.000000m  1.000000 
meas tran maxout max v(net_1) from=0.000000a  to=1.000000 
hardcopy plot1.ps v(net_1) 
hardcopy plot2.ps v(net_3)-v(net_2)


.endc
.end
